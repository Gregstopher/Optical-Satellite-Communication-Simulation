// File: main.sv
// Description: ELEX 7660 main top-level module.
// Author: Taewoo Kim & Greg Kirk
// Date: 2024-04-03
// Last updated: 2024-04-03

module main ( input logic CLOCK_50,       // 50 MHz clock
              output logic [7:0] leds,    // 7-seg LED enables
              output logic [3:0] ct,  // digit cathodes
				  output logic [0:0] GPIO_0,
				  input logic data_input,
              input s1, s2, //pushbuttons		
			     output logic lcd_sda,           // SPI data signal to LCD
				  output logic lcd_scl,           // SPI clock signal to LCD
				  output logic lcd_cs,            // SPI chip select signal to LCD
				  output logic lcd_rs,            // LCD data/command signal
				  output logic lcd_rst,           // LCD reset signal
				  output logic red, green, blue   // RGB LED signals  
            );  
				
				
////////////Soft Processor instantiation////////////////////////////////////////////

    // gpio signal from processor PIN ASSIGNMNET unknown rn
    //logic [7:0] gpio;  

    // instantiate processor system
    soft_processor u0 (
		.clk_clk             (CLOCK_50),//MATCHED
		.gpio_export         (pattern),//MODIFY THIS TO TAKE THE VALUE READ FROM THE LASER
		.reset_reset_n       (s1),
		.spi_0_external_MISO ('0),//unused
		.spi_0_external_MOSI (lcd_sda),//unused
		.spi_0_external_SCLK (lcd_scl),//unused
		.spi_0_external_SS_n (lcd_cs)//unused
	);
 	
    // control the display data/command (lcd_rs) with gpio[0] from processor UNUSED
    //assign lcd_rs = gpio[0];
	
    // control active low display reset (lcd_rst) with gpio[1] from processor UNUSED
    //assign lcd_rst = gpio[1];

	// turn off the RGB LED on the BoosterPack
	assign {red, green, blue} = {'1,'0,'1};
/////////////////////////////////////////////////////////////////////				
				
	
    //7-segment logics
   logic [1:0] digit;           // select digit to display
   logic [3:0] disp_digit;      // current digit of count to display
   logic [15:0] clk_div_count;  // count used to divide clock

   //for freqGen
   logic new_clk;              //secondary clock speed generated by freqgen

   //for sigGen
	
	
   logic [7:0] pattern ;         //Used to send our pattern to sigGen

	
	logic result;                // holds our output from sigGen
	
	logic data_valid;
	logic [7:0] output_data;//data that the laser recieved THIS IS A RECIEVER SIGNAL
   //assign pattern = 
	logic [1:0] pattern_index;  // Goes from 0 to 3
	logic [7:0] current_pattern;
	assign current_pattern = pattern[pattern_index];

	
   // instantiate modules to implement design
   decode2 decode2_0 (.digit, .ct) ;
   decode7 decode7_0 (.num(disp_digit), .leds) ;

   freqgen  #(.FCLK(50000000)) freqgen_0 (.clk(CLOCK_50), .freq(32'd10), .reset_n(s1), .new_freq(new_clk));
   siggen siggen_0 (.pattern(current_pattern),.clk(new_clk), .rst_n(s1), .out_bit(result));
	uart_rx  #(.CLKS_PER_BIT(5208)) uart_rx_0 (.clk(CLOCK_50), .rst_n(s2), .rx_serial(data_input), .data(output_data), .data_valid(data_valid));
	 
	 
	// use count to divide clock and generate a 2 bit digit counter to determine which digit to display
   always_ff @(posedge CLOCK_50) 
     clk_div_count <= clk_div_count + 1'b1 ;

   // assign the top two bits of count to select digit to display
   assign digit = clk_div_count[15:14]; 
	
	assign GPIO_0 = result;
	

  // Select digit to display (disp_digit)
  // Left two digits (3,2) display encoder 1 hex count and right two digits (1,0) display encoder 2 hex count
  always_comb begin
 disp_digit = 4'b0; //assign to 0 on first run
 
	case (digit)
        2'b00: disp_digit = result;  // Encoder 2 Ones place
        2'b01: disp_digit = output_data[3:0];	//output_data[3:0];  // Encoder 2 Tens place
        2'b10: disp_digit = output_data[7:4];  // Encoder 1 Ones place
        2'b11: disp_digit = data_input;  // Encoder 1 Tens place
    endcase  
  end  
  
  logic [25:0] send_timer;
  
  // clock divider to adjust the delay between characters

	

endmodule

