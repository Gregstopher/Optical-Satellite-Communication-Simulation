// File: lab4.sv
// Description: ELEX 7660 lab4 top-level module. uses encoder to choose ADC channel and read from the analog input
// Author: Robert Trost & Greg Kirk (modified)
// Date: 2024-02-05

module main ( input logic CLOCK_50,       // 50 MHz clock
              output logic [7:0] leds,    // 7-seg LED enables
              output logic [3:0] ct,  // digit cathodes
				  output logic [0:0] GPIO_0,
              input s1, s2 //pushbuttons		
            );  //speaker output

    //7-segment logics
   logic [1:0] digit;           // select digit to display
   logic [3:0] disp_digit;      // current digit of count to display
   logic [15:0] clk_div_count;  // count used to divide clock

   //for freqGen
   logic new_clk;              //secondary clock speed generated by freqgen

   //for sigGen
   logic [6:0] pattern;         //Used to send our pattern to sigGen
   logic result;                // holds our output from sigGen

   assign pattern = 7'b1001010;
   
   // instantiate modules to implement design
   decode2 decode2_0 (.digit, .ct) ;
   decode7 decode7_0 (.num(disp_digit), .leds) ;

   freqgen  #(.FCLK(50000000)) freqgen_0 (.clk(CLOCK_50), .freq(32'd2000, .reset_n(s1), .new_freq(new_clk));
   siggen siggen_0 (.pattern(pattern),.clk(new_clk), .rst_n(s1),.out_bit(result));
   

   // use count to divide clock and generate a 2 bit digit counter to determine which digit to display
   always_ff @(posedge CLOCK_50) 
     clk_div_count <= clk_div_count + 1'b1 ;

   // assign the top two bits of count to select digit to display
   assign digit = clk_div_count[15:14]; 
	
	assign GPIO_0 = result;
	

  // Select digit to display (disp_digit)
  // Left two digits (3,2) display encoder 1 hex count and right two digits (1,0) display encoder 2 hex count
  always_comb begin
 disp_digit = 4'b0; //assign to 0 on first run
 
case (digit)
        2'b00: disp_digit = result;  // Encoder 2 Ones place
        2'b01: disp_digit = 4'b0;  // Encoder 2 Tens place
        2'b10: disp_digit = 4'b0;  // Encoder 1 Ones place
        2'b11: disp_digit = 4'b0;  // Encoder 1 Tens place
    endcase  
  end  

endmodule

